// Copyright 2006, 2007 Dennis van Weeren
//
// This file is part of Minimig
//
// Minimig is free software; you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation; either version 3 of the License, or
// (at your option) any later version.
//
// Minimig is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>.
//
//
//
// This is the Minimig boot rom
// The bootrom contains code for early startup of the Minimig.
// The bootrom will download the kickstart rom image trough the floppy 
// interface to the kickstart ram area. 
//
// 11-04-2005	-removed rd signal because it is no longer necessary
// 19-04-2005	-expanded to 2Kbyte address space
// 21-12-2005	-added rd input
// 27-11-2006	-rom now implemented using blockram

module bootrom(clk,aen,rd,address,dataout);
input 	clk;					//bus clock
input 	aen;    				//rom enable
input	rd;					//bus read
input 	[10:1]address;			//address in
output 	[15:0]dataout;	 		//data out

reg 		[15:0]dataout;
reg	 	[10:1]romaddress;
reg		[15:0]romdata;

//use clocked address to infer blockram
always @(negedge clk)
	romaddress[10:1]<=address[10:1];

//the rom itself
//if all goes well this rom will be implemented using blockram
always @(romaddress)
begin	
	case(romaddress)
		0000:	romdata[15:0]=16'h0007;
		0001:	romdata[15:0]=16'h0100;
		0002:	romdata[15:0]=16'h0000;
		0003:	romdata[15:0]=16'h0100;
		0004:	romdata[15:0]=16'h0000;
		0005:	romdata[15:0]=16'h0000;
		0006:	romdata[15:0]=16'h0000;
		0007:	romdata[15:0]=16'h0000;
		0008:	romdata[15:0]=16'h0000;
		0009:	romdata[15:0]=16'h0000;
		0010:	romdata[15:0]=16'h0000;
		0011:	romdata[15:0]=16'h0000;
		0012:	romdata[15:0]=16'h0000;
		0013:	romdata[15:0]=16'h0000;
		0014:	romdata[15:0]=16'h0000;
		0015:	romdata[15:0]=16'h0000;
		0016:	romdata[15:0]=16'h0000;
		0017:	romdata[15:0]=16'h0000;
		0018:	romdata[15:0]=16'h0000;
		0019:	romdata[15:0]=16'h0000;
		0020:	romdata[15:0]=16'h0000;
		0021:	romdata[15:0]=16'h0000;
		0022:	romdata[15:0]=16'h0000;
		0023:	romdata[15:0]=16'h0000;
		0024:	romdata[15:0]=16'h0000;
		0025:	romdata[15:0]=16'h0000;
		0026:	romdata[15:0]=16'h0000;
		0027:	romdata[15:0]=16'h0000;
		0028:	romdata[15:0]=16'h0000;
		0029:	romdata[15:0]=16'h0000;
		0030:	romdata[15:0]=16'h0000;
		0031:	romdata[15:0]=16'h0000;
		0032:	romdata[15:0]=16'h0000;
		0033:	romdata[15:0]=16'h0000;
		0034:	romdata[15:0]=16'h0000;
		0035:	romdata[15:0]=16'h0000;
		0036:	romdata[15:0]=16'h0000;
		0037:	romdata[15:0]=16'h0000;
		0038:	romdata[15:0]=16'h0000;
		0039:	romdata[15:0]=16'h0000;
		0040:	romdata[15:0]=16'h0000;
		0041:	romdata[15:0]=16'h0000;
		0042:	romdata[15:0]=16'h0000;
		0043:	romdata[15:0]=16'h0000;
		0044:	romdata[15:0]=16'h0000;
		0045:	romdata[15:0]=16'h0000;
		0046:	romdata[15:0]=16'h0000;
		0047:	romdata[15:0]=16'h0000;
		0048:	romdata[15:0]=16'h0000;
		0049:	romdata[15:0]=16'h0000;
		0050:	romdata[15:0]=16'h0000;
		0051:	romdata[15:0]=16'h0000;
		0052:	romdata[15:0]=16'h0000;
		0053:	romdata[15:0]=16'h0000;
		0054:	romdata[15:0]=16'h0000;
		0055:	romdata[15:0]=16'h0000;
		0056:	romdata[15:0]=16'h0000;
		0057:	romdata[15:0]=16'h0000;
		0058:	romdata[15:0]=16'h0000;
		0059:	romdata[15:0]=16'h0000;
		0060:	romdata[15:0]=16'h0000;
		0061:	romdata[15:0]=16'h0000;
		0062:	romdata[15:0]=16'h0000;
		0063:	romdata[15:0]=16'h0000;
		0064:	romdata[15:0]=16'h0000;
		0065:	romdata[15:0]=16'h0000;
		0066:	romdata[15:0]=16'h0000;
		0067:	romdata[15:0]=16'h0000;
		0068:	romdata[15:0]=16'h0000;
		0069:	romdata[15:0]=16'h0000;
		0070:	romdata[15:0]=16'h0000;
		0071:	romdata[15:0]=16'h0000;
		0072:	romdata[15:0]=16'h0000;
		0073:	romdata[15:0]=16'h0000;
		0074:	romdata[15:0]=16'h0000;
		0075:	romdata[15:0]=16'h0000;
		0076:	romdata[15:0]=16'h0000;
		0077:	romdata[15:0]=16'h0000;
		0078:	romdata[15:0]=16'h0000;
		0079:	romdata[15:0]=16'h0000;
		0080:	romdata[15:0]=16'h0000;
		0081:	romdata[15:0]=16'h0000;
		0082:	romdata[15:0]=16'h0000;
		0083:	romdata[15:0]=16'h0000;
		0084:	romdata[15:0]=16'h0000;
		0085:	romdata[15:0]=16'h0000;
		0086:	romdata[15:0]=16'h0000;
		0087:	romdata[15:0]=16'h0000;
		0088:	romdata[15:0]=16'h0000;
		0089:	romdata[15:0]=16'h0000;
		0090:	romdata[15:0]=16'h0000;
		0091:	romdata[15:0]=16'h0000;
		0092:	romdata[15:0]=16'h0000;
		0093:	romdata[15:0]=16'h0000;
		0094:	romdata[15:0]=16'h0000;
		0095:	romdata[15:0]=16'h0000;
		0096:	romdata[15:0]=16'h0000;
		0097:	romdata[15:0]=16'h0000;
		0098:	romdata[15:0]=16'h0000;
		0099:	romdata[15:0]=16'h0000;
		0100:	romdata[15:0]=16'h0000;
		0101:	romdata[15:0]=16'h0000;
		0102:	romdata[15:0]=16'h0000;
		0103:	romdata[15:0]=16'h0000;
		0104:	romdata[15:0]=16'h0000;
		0105:	romdata[15:0]=16'h0000;
		0106:	romdata[15:0]=16'h0000;
		0107:	romdata[15:0]=16'h0000;
		0108:	romdata[15:0]=16'h0000;
		0109:	romdata[15:0]=16'h0000;
		0110:	romdata[15:0]=16'h0000;
		0111:	romdata[15:0]=16'h0000;
		0112:	romdata[15:0]=16'h0000;
		0113:	romdata[15:0]=16'h0000;
		0114:	romdata[15:0]=16'h0000;
		0115:	romdata[15:0]=16'h0000;
		0116:	romdata[15:0]=16'h0000;
		0117:	romdata[15:0]=16'h0000;
		0118:	romdata[15:0]=16'h0000;
		0119:	romdata[15:0]=16'h0000;
		0120:	romdata[15:0]=16'h0000;
		0121:	romdata[15:0]=16'h0000;
		0122:	romdata[15:0]=16'h0000;
		0123:	romdata[15:0]=16'h0000;
		0124:	romdata[15:0]=16'h0000;
		0125:	romdata[15:0]=16'h0000;
		0126:	romdata[15:0]=16'h0000;
		0127:	romdata[15:0]=16'h0000;
		0128:	romdata[15:0]=16'h41F9;
		0129:	romdata[15:0]=16'h00DF;
		0130:	romdata[15:0]=16'hF000;
		0131:	romdata[15:0]=16'h43F9;
		0132:	romdata[15:0]=16'h00BF;
		0133:	romdata[15:0]=16'hE001;
		0134:	romdata[15:0]=16'h45F9;
		0135:	romdata[15:0]=16'h00BF;
		0136:	romdata[15:0]=16'hD000;
		0137:	romdata[15:0]=16'h47F9;
		0138:	romdata[15:0]=16'h00F8;
		0139:	romdata[15:0]=16'h0000;
		0140:	romdata[15:0]=16'h157C;
		0141:	romdata[15:0]=16'h00F7;
		0142:	romdata[15:0]=16'h0100;
		0143:	romdata[15:0]=16'h157C;
		0144:	romdata[15:0]=16'h00FF;
		0145:	romdata[15:0]=16'h0300;
		0146:	romdata[15:0]=16'h317C;
		0147:	romdata[15:0]=16'h001E;
		0148:	romdata[15:0]=16'h0032;
		0149:	romdata[15:0]=16'h317C;
		0150:	romdata[15:0]=16'h7000;
		0151:	romdata[15:0]=16'h009A;
		0152:	romdata[15:0]=16'h317C;
		0153:	romdata[15:0]=16'h7FFF;
		0154:	romdata[15:0]=16'h009C;
		0155:	romdata[15:0]=16'h317C;
		0156:	romdata[15:0]=16'h8210;
		0157:	romdata[15:0]=16'h0096;
		0158:	romdata[15:0]=16'h317C;
		0159:	romdata[15:0]=16'h7FFF;
		0160:	romdata[15:0]=16'h009E;
		0161:	romdata[15:0]=16'h6100;
		0162:	romdata[15:0]=16'h0028;
		0163:	romdata[15:0]=16'h08AA;
		0164:	romdata[15:0]=16'h0001;
		0165:	romdata[15:0]=16'h0100;
		0166:	romdata[15:0]=16'h6100;
		0167:	romdata[15:0]=16'h003A;
		0168:	romdata[15:0]=16'h6100;
		0169:	romdata[15:0]=16'h0062;
		0170:	romdata[15:0]=16'hB7FC;
		0171:	romdata[15:0]=16'h0100;
		0172:	romdata[15:0]=16'h0000;
		0173:	romdata[15:0]=16'h6700;
		0174:	romdata[15:0]=16'h0070;
		0175:	romdata[15:0]=16'h08AA;
		0176:	romdata[15:0]=16'h0000;
		0177:	romdata[15:0]=16'h0100;
		0178:	romdata[15:0]=16'h08EA;
		0179:	romdata[15:0]=16'h0000;
		0180:	romdata[15:0]=16'h0100;
		0181:	romdata[15:0]=16'h60E0;
		0182:	romdata[15:0]=16'h103C;
		0183:	romdata[15:0]=16'h00FF;
		0184:	romdata[15:0]=16'h08EA;
		0185:	romdata[15:0]=16'h0001;
		0186:	romdata[15:0]=16'h0100;
		0187:	romdata[15:0]=16'h08AA;
		0188:	romdata[15:0]=16'h0000;
		0189:	romdata[15:0]=16'h0100;
		0190:	romdata[15:0]=16'h08EA;
		0191:	romdata[15:0]=16'h0000;
		0192:	romdata[15:0]=16'h0100;
		0193:	romdata[15:0]=16'h51C8;
		0194:	romdata[15:0]=16'hFFF2;
		0195:	romdata[15:0]=16'h4E75;
		0196:	romdata[15:0]=16'h217C;
		0197:	romdata[15:0]=16'h0001;
		0198:	romdata[15:0]=16'h0000;
		0199:	romdata[15:0]=16'h0020;
		0200:	romdata[15:0]=16'h317C;
		0201:	romdata[15:0]=16'h0002;
		0202:	romdata[15:0]=16'h009C;
		0203:	romdata[15:0]=16'h317C;
		0204:	romdata[15:0]=16'hA000;
		0205:	romdata[15:0]=16'h0024;
		0206:	romdata[15:0]=16'h317C;
		0207:	romdata[15:0]=16'hA000;
		0208:	romdata[15:0]=16'h0024;
		0209:	romdata[15:0]=16'h3028;
		0210:	romdata[15:0]=16'h001E;
		0211:	romdata[15:0]=16'hC07C;
		0212:	romdata[15:0]=16'h0002;
		0213:	romdata[15:0]=16'h67F6;
		0214:	romdata[15:0]=16'h317C;
		0215:	romdata[15:0]=16'h4000;
		0216:	romdata[15:0]=16'h0024;
		0217:	romdata[15:0]=16'h4E75;
		0218:	romdata[15:0]=16'h303C;
		0219:	romdata[15:0]=16'h0FFF;
		0220:	romdata[15:0]=16'h49F9;
		0221:	romdata[15:0]=16'h0001;
		0222:	romdata[15:0]=16'h0000;
		0223:	romdata[15:0]=16'h221C;
		0224:	romdata[15:0]=16'h26C1;
		0225:	romdata[15:0]=16'h3141;
		0226:	romdata[15:0]=16'h0180;
		0227:	romdata[15:0]=16'h51C8;
		0228:	romdata[15:0]=16'hFFF6;
		0229:	romdata[15:0]=16'h4E75;
		0230:	romdata[15:0]=16'h13C0;
		0231:	romdata[15:0]=16'h00BF;
		0232:	romdata[15:0]=16'hC000;
		0233:	romdata[15:0]=16'h60F8;
		0234:	romdata[15:0]=16'h0000;
		0235:	romdata[15:0]=16'h0000;
		0236:	romdata[15:0]=16'h0000;
		0237:	romdata[15:0]=16'h0000;
		0238:	romdata[15:0]=16'h0000;
		0239:	romdata[15:0]=16'h0000;
		0240:	romdata[15:0]=16'h0000;
		0241:	romdata[15:0]=16'h0000;
		0242:	romdata[15:0]=16'h0000;
		0243:	romdata[15:0]=16'h0000;
		0244:	romdata[15:0]=16'h0000;
		0245:	romdata[15:0]=16'h0000;
		0246:	romdata[15:0]=16'h0000;
		0247:	romdata[15:0]=16'h0000;
		0248:	romdata[15:0]=16'h0000;
		0249:	romdata[15:0]=16'h0000;
		0250:	romdata[15:0]=16'h0000;
		0251:	romdata[15:0]=16'h0000;
		0252:	romdata[15:0]=16'h0000;
		0253:	romdata[15:0]=16'h0000;
		0254:	romdata[15:0]=16'h0000;
		0255:	romdata[15:0]=16'h0000;
		0256:	romdata[15:0]=16'h0000;
		0257:	romdata[15:0]=16'h0000;
		0258:	romdata[15:0]=16'h0000;
		0259:	romdata[15:0]=16'h0000;
		0260:	romdata[15:0]=16'h0000;
		0261:	romdata[15:0]=16'h0000;
		0262:	romdata[15:0]=16'h0000;
		0263:	romdata[15:0]=16'h0000;
		0264:	romdata[15:0]=16'h0000;
		0265:	romdata[15:0]=16'h0000;
		0266:	romdata[15:0]=16'h0000;
		0267:	romdata[15:0]=16'h0000;
		0268:	romdata[15:0]=16'h0000;
		0269:	romdata[15:0]=16'h0000;
		0270:	romdata[15:0]=16'h0000;
		0271:	romdata[15:0]=16'h0000;
		0272:	romdata[15:0]=16'h0000;
		0273:	romdata[15:0]=16'h0000;
		0274:	romdata[15:0]=16'h0000;
		0275:	romdata[15:0]=16'h0000;
		0276:	romdata[15:0]=16'h0000;
		0277:	romdata[15:0]=16'h0000;
		0278:	romdata[15:0]=16'h0000;
		0279:	romdata[15:0]=16'h0000;
		0280:	romdata[15:0]=16'h0000;
		0281:	romdata[15:0]=16'h0000;
		0282:	romdata[15:0]=16'h0000;
		0283:	romdata[15:0]=16'h0000;
		0284:	romdata[15:0]=16'h0000;
		0285:	romdata[15:0]=16'h0000;
		0286:	romdata[15:0]=16'h0000;
		0287:	romdata[15:0]=16'h0000;
		0288:	romdata[15:0]=16'h0000;
		0289:	romdata[15:0]=16'h0000;
		0290:	romdata[15:0]=16'h0000;
		0291:	romdata[15:0]=16'h0000;
		0292:	romdata[15:0]=16'h0000;
		0293:	romdata[15:0]=16'h0000;
		0294:	romdata[15:0]=16'h0000;
		0295:	romdata[15:0]=16'h0000;
		0296:	romdata[15:0]=16'h0000;
		0297:	romdata[15:0]=16'h0000;
		0298:	romdata[15:0]=16'h0000;
		0299:	romdata[15:0]=16'h0000;
		0300:	romdata[15:0]=16'h0000;
		0301:	romdata[15:0]=16'h0000;
		0302:	romdata[15:0]=16'h0000;
		0303:	romdata[15:0]=16'h0000;
		0304:	romdata[15:0]=16'h0000;
		0305:	romdata[15:0]=16'h0000;
		0306:	romdata[15:0]=16'h0000;
		0307:	romdata[15:0]=16'h0000;
		0308:	romdata[15:0]=16'h0000;
		0309:	romdata[15:0]=16'h0000;
		0310:	romdata[15:0]=16'h0000;
		0311:	romdata[15:0]=16'h0000;
		0312:	romdata[15:0]=16'h0000;
		0313:	romdata[15:0]=16'h0000;
		0314:	romdata[15:0]=16'h0000;
		0315:	romdata[15:0]=16'h0000;
		0316:	romdata[15:0]=16'h0000;
		0317:	romdata[15:0]=16'h0000;
		0318:	romdata[15:0]=16'h0000;
		0319:	romdata[15:0]=16'h0000;
		0320:	romdata[15:0]=16'h0000;
		0321:	romdata[15:0]=16'h0000;
		0322:	romdata[15:0]=16'h0000;
		0323:	romdata[15:0]=16'h0000;
		0324:	romdata[15:0]=16'h0000;
		0325:	romdata[15:0]=16'h0000;
		0326:	romdata[15:0]=16'h0000;
		0327:	romdata[15:0]=16'h0000;
		0328:	romdata[15:0]=16'h0000;
		0329:	romdata[15:0]=16'h0000;
		0330:	romdata[15:0]=16'h0000;
		0331:	romdata[15:0]=16'h0000;
		0332:	romdata[15:0]=16'h0000;
		0333:	romdata[15:0]=16'h0000;
		0334:	romdata[15:0]=16'h0000;
		0335:	romdata[15:0]=16'h0000;
		0336:	romdata[15:0]=16'h0000;
		0337:	romdata[15:0]=16'h0000;
		0338:	romdata[15:0]=16'h0000;
		0339:	romdata[15:0]=16'h0000;
		0340:	romdata[15:0]=16'h0000;
		0341:	romdata[15:0]=16'h0000;
		0342:	romdata[15:0]=16'h0000;
		0343:	romdata[15:0]=16'h0000;
		0344:	romdata[15:0]=16'h0000;
		0345:	romdata[15:0]=16'h0000;
		0346:	romdata[15:0]=16'h0000;
		0347:	romdata[15:0]=16'h0000;
		0348:	romdata[15:0]=16'h0000;
		0349:	romdata[15:0]=16'h0000;
		0350:	romdata[15:0]=16'h0000;
		0351:	romdata[15:0]=16'h0000;
		0352:	romdata[15:0]=16'h0000;
		0353:	romdata[15:0]=16'h0000;
		0354:	romdata[15:0]=16'h0000;
		0355:	romdata[15:0]=16'h0000;
		0356:	romdata[15:0]=16'h0000;
		0357:	romdata[15:0]=16'h0000;
		0358:	romdata[15:0]=16'h0000;
		0359:	romdata[15:0]=16'h0000;
		0360:	romdata[15:0]=16'h0000;
		0361:	romdata[15:0]=16'h0000;
		0362:	romdata[15:0]=16'h0000;
		0363:	romdata[15:0]=16'h0000;
		0364:	romdata[15:0]=16'h0000;
		0365:	romdata[15:0]=16'h0000;
		0366:	romdata[15:0]=16'h0000;
		0367:	romdata[15:0]=16'h0000;
		0368:	romdata[15:0]=16'h0000;
		0369:	romdata[15:0]=16'h0000;
		0370:	romdata[15:0]=16'h0000;
		0371:	romdata[15:0]=16'h0000;
		0372:	romdata[15:0]=16'h0000;
		0373:	romdata[15:0]=16'h0000;
		0374:	romdata[15:0]=16'h0000;
		0375:	romdata[15:0]=16'h0000;
		0376:	romdata[15:0]=16'h0000;
		0377:	romdata[15:0]=16'h0000;
		0378:	romdata[15:0]=16'h0000;
		0379:	romdata[15:0]=16'h0000;
		0380:	romdata[15:0]=16'h0000;
		0381:	romdata[15:0]=16'h0000;
		0382:	romdata[15:0]=16'h0000;
		0383:	romdata[15:0]=16'h0000;
		0384:	romdata[15:0]=16'h0000;
		0385:	romdata[15:0]=16'h0000;
		0386:	romdata[15:0]=16'h0000;
		0387:	romdata[15:0]=16'h0000;
		0388:	romdata[15:0]=16'h0000;
		0389:	romdata[15:0]=16'h0000;
		0390:	romdata[15:0]=16'h0000;
		0391:	romdata[15:0]=16'h0000;
		0392:	romdata[15:0]=16'h0000;
		0393:	romdata[15:0]=16'h0000;
		0394:	romdata[15:0]=16'h0000;
		0395:	romdata[15:0]=16'h0000;
		0396:	romdata[15:0]=16'h0000;
		0397:	romdata[15:0]=16'h0000;
		0398:	romdata[15:0]=16'h0000;
		0399:	romdata[15:0]=16'h0000;
		0400:	romdata[15:0]=16'h0000;
		0401:	romdata[15:0]=16'h0000;
		0402:	romdata[15:0]=16'h0000;
		0403:	romdata[15:0]=16'h0000;
		0404:	romdata[15:0]=16'h0000;
		0405:	romdata[15:0]=16'h0000;
		0406:	romdata[15:0]=16'h0000;
		0407:	romdata[15:0]=16'h0000;
		0408:	romdata[15:0]=16'h0000;
		0409:	romdata[15:0]=16'h0000;
		0410:	romdata[15:0]=16'h0000;
		0411:	romdata[15:0]=16'h0000;
		0412:	romdata[15:0]=16'h0000;
		0413:	romdata[15:0]=16'h0000;
		0414:	romdata[15:0]=16'h0000;
		0415:	romdata[15:0]=16'h0000;
		0416:	romdata[15:0]=16'h0000;
		0417:	romdata[15:0]=16'h0000;
		0418:	romdata[15:0]=16'h0000;
		0419:	romdata[15:0]=16'h0000;
		0420:	romdata[15:0]=16'h0000;
		0421:	romdata[15:0]=16'h0000;
		0422:	romdata[15:0]=16'h0000;
		0423:	romdata[15:0]=16'h0000;
		0424:	romdata[15:0]=16'h0000;
		0425:	romdata[15:0]=16'h0000;
		0426:	romdata[15:0]=16'h0000;
		0427:	romdata[15:0]=16'h0000;
		0428:	romdata[15:0]=16'h0000;
		0429:	romdata[15:0]=16'h0000;
		0430:	romdata[15:0]=16'h0000;
		0431:	romdata[15:0]=16'h0000;
		0432:	romdata[15:0]=16'h0000;
		0433:	romdata[15:0]=16'h0000;
		0434:	romdata[15:0]=16'h0000;
		0435:	romdata[15:0]=16'h0000;
		0436:	romdata[15:0]=16'h0000;
		0437:	romdata[15:0]=16'h0000;
		0438:	romdata[15:0]=16'h0000;
		0439:	romdata[15:0]=16'h0000;
		0440:	romdata[15:0]=16'h0000;
		0441:	romdata[15:0]=16'h0000;
		0442:	romdata[15:0]=16'h0000;
		0443:	romdata[15:0]=16'h0000;
		0444:	romdata[15:0]=16'h0000;
		0445:	romdata[15:0]=16'h0000;
		0446:	romdata[15:0]=16'h0000;
		0447:	romdata[15:0]=16'h0000;
		0448:	romdata[15:0]=16'h0000;
		0449:	romdata[15:0]=16'h0000;
		0450:	romdata[15:0]=16'h0000;
		0451:	romdata[15:0]=16'h0000;
		0452:	romdata[15:0]=16'h0000;
		0453:	romdata[15:0]=16'h0000;
		0454:	romdata[15:0]=16'h0000;
		0455:	romdata[15:0]=16'h0000;
		0456:	romdata[15:0]=16'h0000;
		0457:	romdata[15:0]=16'h0000;
		0458:	romdata[15:0]=16'h0000;
		0459:	romdata[15:0]=16'h0000;
		0460:	romdata[15:0]=16'h0000;
		0461:	romdata[15:0]=16'h0000;
		0462:	romdata[15:0]=16'h0000;
		0463:	romdata[15:0]=16'h0000;
		0464:	romdata[15:0]=16'h0000;
		0465:	romdata[15:0]=16'h0000;
		0466:	romdata[15:0]=16'h0000;
		0467:	romdata[15:0]=16'h0000;
		0468:	romdata[15:0]=16'h0000;
		0469:	romdata[15:0]=16'h0000;
		0470:	romdata[15:0]=16'h0000;
		0471:	romdata[15:0]=16'h0000;
		0472:	romdata[15:0]=16'h0000;
		0473:	romdata[15:0]=16'h0000;
		0474:	romdata[15:0]=16'h0000;
		0475:	romdata[15:0]=16'h0000;
		0476:	romdata[15:0]=16'h0000;
		0477:	romdata[15:0]=16'h0000;
		0478:	romdata[15:0]=16'h0000;
		0479:	romdata[15:0]=16'h0000;
		0480:	romdata[15:0]=16'h0000;
		0481:	romdata[15:0]=16'h0000;
		0482:	romdata[15:0]=16'h0000;
		0483:	romdata[15:0]=16'h0000;
		0484:	romdata[15:0]=16'h0000;
		0485:	romdata[15:0]=16'h0000;
		0486:	romdata[15:0]=16'h0000;
		0487:	romdata[15:0]=16'h0000;
		0488:	romdata[15:0]=16'h0000;
		0489:	romdata[15:0]=16'h0000;
		0490:	romdata[15:0]=16'h0000;
		0491:	romdata[15:0]=16'h0000;
		0492:	romdata[15:0]=16'h0000;
		0493:	romdata[15:0]=16'h0000;
		0494:	romdata[15:0]=16'h0000;
		0495:	romdata[15:0]=16'h0000;
		0496:	romdata[15:0]=16'h0000;
		0497:	romdata[15:0]=16'h0000;
		0498:	romdata[15:0]=16'h0000;
		0499:	romdata[15:0]=16'h0000;
		0500:	romdata[15:0]=16'h0000;
		0501:	romdata[15:0]=16'h0000;
		0502:	romdata[15:0]=16'h0000;
		0503:	romdata[15:0]=16'h0000;
		0504:	romdata[15:0]=16'h0000;
		0505:	romdata[15:0]=16'h0000;
		0506:	romdata[15:0]=16'h0000;
		0507:	romdata[15:0]=16'h0000;
		0508:	romdata[15:0]=16'h0000;
		0509:	romdata[15:0]=16'h0000;
		0510:	romdata[15:0]=16'h0000;
		0511:	romdata[15:0]=16'h0000;
		0512:	romdata[15:0]=16'h0000;
		0513:	romdata[15:0]=16'h0000;
		0514:	romdata[15:0]=16'h0000;
		0515:	romdata[15:0]=16'h0000;
		0516:	romdata[15:0]=16'h0000;
		0517:	romdata[15:0]=16'h0000;
		0518:	romdata[15:0]=16'h0000;
		0519:	romdata[15:0]=16'h0000;
		0520:	romdata[15:0]=16'h0000;
		0521:	romdata[15:0]=16'h0000;
		0522:	romdata[15:0]=16'h0000;
		0523:	romdata[15:0]=16'h0000;
		0524:	romdata[15:0]=16'h0000;
		0525:	romdata[15:0]=16'h0000;
		0526:	romdata[15:0]=16'h0000;
		0527:	romdata[15:0]=16'h0000;
		0528:	romdata[15:0]=16'h0000;
		0529:	romdata[15:0]=16'h0000;
		0530:	romdata[15:0]=16'h0000;
		0531:	romdata[15:0]=16'h0000;
		0532:	romdata[15:0]=16'h0000;
		0533:	romdata[15:0]=16'h0000;
		0534:	romdata[15:0]=16'h0000;
		0535:	romdata[15:0]=16'h0000;
		0536:	romdata[15:0]=16'h0000;
		0537:	romdata[15:0]=16'h0000;
		0538:	romdata[15:0]=16'h0000;
		0539:	romdata[15:0]=16'h0000;
		0540:	romdata[15:0]=16'h0000;
		0541:	romdata[15:0]=16'h0000;
		0542:	romdata[15:0]=16'h0000;
		0543:	romdata[15:0]=16'h0000;
		0544:	romdata[15:0]=16'h0000;
		0545:	romdata[15:0]=16'h0000;
		0546:	romdata[15:0]=16'h0000;
		0547:	romdata[15:0]=16'h0000;
		0548:	romdata[15:0]=16'h0000;
		0549:	romdata[15:0]=16'h0000;
		0550:	romdata[15:0]=16'h0000;
		0551:	romdata[15:0]=16'h0000;
		0552:	romdata[15:0]=16'h0000;
		0553:	romdata[15:0]=16'h0000;
		0554:	romdata[15:0]=16'h0000;
		0555:	romdata[15:0]=16'h0000;
		0556:	romdata[15:0]=16'h0000;
		0557:	romdata[15:0]=16'h0000;
		0558:	romdata[15:0]=16'h0000;
		0559:	romdata[15:0]=16'h0000;
		0560:	romdata[15:0]=16'h0000;
		0561:	romdata[15:0]=16'h0000;
		0562:	romdata[15:0]=16'h0000;
		0563:	romdata[15:0]=16'h0000;
		0564:	romdata[15:0]=16'h0000;
		0565:	romdata[15:0]=16'h0000;
		0566:	romdata[15:0]=16'h0000;
		0567:	romdata[15:0]=16'h0000;
		0568:	romdata[15:0]=16'h0000;
		0569:	romdata[15:0]=16'h0000;
		0570:	romdata[15:0]=16'h0000;
		0571:	romdata[15:0]=16'h0000;
		0572:	romdata[15:0]=16'h0000;
		0573:	romdata[15:0]=16'h0000;
		0574:	romdata[15:0]=16'h0000;
		0575:	romdata[15:0]=16'h0000;
		0576:	romdata[15:0]=16'h0000;
		0577:	romdata[15:0]=16'h0000;
		0578:	romdata[15:0]=16'h0000;
		0579:	romdata[15:0]=16'h0000;
		0580:	romdata[15:0]=16'h0000;
		0581:	romdata[15:0]=16'h0000;
		0582:	romdata[15:0]=16'h0000;
		0583:	romdata[15:0]=16'h0000;
		0584:	romdata[15:0]=16'h0000;
		0585:	romdata[15:0]=16'h0000;
		0586:	romdata[15:0]=16'h0000;
		0587:	romdata[15:0]=16'h0000;
		0588:	romdata[15:0]=16'h0000;
		0589:	romdata[15:0]=16'h0000;
		0590:	romdata[15:0]=16'h0000;
		0591:	romdata[15:0]=16'h0000;
		0592:	romdata[15:0]=16'h0000;
		0593:	romdata[15:0]=16'h0000;
		0594:	romdata[15:0]=16'h0000;
		0595:	romdata[15:0]=16'h0000;
		0596:	romdata[15:0]=16'h0000;
		0597:	romdata[15:0]=16'h0000;
		0598:	romdata[15:0]=16'h0000;
		0599:	romdata[15:0]=16'h0000;
		0600:	romdata[15:0]=16'h0000;
		0601:	romdata[15:0]=16'h0000;
		0602:	romdata[15:0]=16'h0000;
		0603:	romdata[15:0]=16'h0000;
		0604:	romdata[15:0]=16'h0000;
		0605:	romdata[15:0]=16'h0000;
		0606:	romdata[15:0]=16'h0000;
		0607:	romdata[15:0]=16'h0000;
		0608:	romdata[15:0]=16'h0000;
		0609:	romdata[15:0]=16'h0000;
		0610:	romdata[15:0]=16'h0000;
		0611:	romdata[15:0]=16'h0000;
		0612:	romdata[15:0]=16'h0000;
		0613:	romdata[15:0]=16'h0000;
		0614:	romdata[15:0]=16'h0000;
		0615:	romdata[15:0]=16'h0000;
		0616:	romdata[15:0]=16'h0000;
		0617:	romdata[15:0]=16'h0000;
		0618:	romdata[15:0]=16'h0000;
		0619:	romdata[15:0]=16'h0000;
		0620:	romdata[15:0]=16'h0000;
		0621:	romdata[15:0]=16'h0000;
		0622:	romdata[15:0]=16'h0000;
		0623:	romdata[15:0]=16'h0000;
		0624:	romdata[15:0]=16'h0000;
		0625:	romdata[15:0]=16'h0000;
		0626:	romdata[15:0]=16'h0000;
		0627:	romdata[15:0]=16'h0000;
		0628:	romdata[15:0]=16'h0000;
		0629:	romdata[15:0]=16'h0000;
		0630:	romdata[15:0]=16'h0000;
		0631:	romdata[15:0]=16'h0000;
		0632:	romdata[15:0]=16'h0000;
		0633:	romdata[15:0]=16'h0000;
		0634:	romdata[15:0]=16'h0000;
		0635:	romdata[15:0]=16'h0000;
		0636:	romdata[15:0]=16'h0000;
		0637:	romdata[15:0]=16'h0000;
		0638:	romdata[15:0]=16'h0000;
		0639:	romdata[15:0]=16'h0000;
		0640:	romdata[15:0]=16'h0000;
		0641:	romdata[15:0]=16'h0000;
		0642:	romdata[15:0]=16'h0000;
		0643:	romdata[15:0]=16'h0000;
		0644:	romdata[15:0]=16'h0000;
		0645:	romdata[15:0]=16'h0000;
		0646:	romdata[15:0]=16'h0000;
		0647:	romdata[15:0]=16'h0000;
		0648:	romdata[15:0]=16'h0000;
		0649:	romdata[15:0]=16'h0000;
		0650:	romdata[15:0]=16'h0000;
		0651:	romdata[15:0]=16'h0000;
		0652:	romdata[15:0]=16'h0000;
		0653:	romdata[15:0]=16'h0000;
		0654:	romdata[15:0]=16'h0000;
		0655:	romdata[15:0]=16'h0000;
		0656:	romdata[15:0]=16'h0000;
		0657:	romdata[15:0]=16'h0000;
		0658:	romdata[15:0]=16'h0000;
		0659:	romdata[15:0]=16'h0000;
		0660:	romdata[15:0]=16'h0000;
		0661:	romdata[15:0]=16'h0000;
		0662:	romdata[15:0]=16'h0000;
		0663:	romdata[15:0]=16'h0000;
		0664:	romdata[15:0]=16'h0000;
		0665:	romdata[15:0]=16'h0000;
		0666:	romdata[15:0]=16'h0000;
		0667:	romdata[15:0]=16'h0000;
		0668:	romdata[15:0]=16'h0000;
		0669:	romdata[15:0]=16'h0000;
		0670:	romdata[15:0]=16'h0000;
		0671:	romdata[15:0]=16'h0000;
		0672:	romdata[15:0]=16'h0000;
		0673:	romdata[15:0]=16'h0000;
		0674:	romdata[15:0]=16'h0000;
		0675:	romdata[15:0]=16'h0000;
		0676:	romdata[15:0]=16'h0000;
		0677:	romdata[15:0]=16'h0000;
		0678:	romdata[15:0]=16'h0000;
		0679:	romdata[15:0]=16'h0000;
		0680:	romdata[15:0]=16'h0000;
		0681:	romdata[15:0]=16'h0000;
		0682:	romdata[15:0]=16'h0000;
		0683:	romdata[15:0]=16'h0000;
		0684:	romdata[15:0]=16'h0000;
		0685:	romdata[15:0]=16'h0000;
		0686:	romdata[15:0]=16'h0000;
		0687:	romdata[15:0]=16'h0000;
		0688:	romdata[15:0]=16'h0000;
		0689:	romdata[15:0]=16'h0000;
		0690:	romdata[15:0]=16'h0000;
		0691:	romdata[15:0]=16'h0000;
		0692:	romdata[15:0]=16'h0000;
		0693:	romdata[15:0]=16'h0000;
		0694:	romdata[15:0]=16'h0000;
		0695:	romdata[15:0]=16'h0000;
		0696:	romdata[15:0]=16'h0000;
		0697:	romdata[15:0]=16'h0000;
		0698:	romdata[15:0]=16'h0000;
		0699:	romdata[15:0]=16'h0000;
		0700:	romdata[15:0]=16'h0000;
		0701:	romdata[15:0]=16'h0000;
		0702:	romdata[15:0]=16'h0000;
		0703:	romdata[15:0]=16'h0000;
		0704:	romdata[15:0]=16'h0000;
		0705:	romdata[15:0]=16'h0000;
		0706:	romdata[15:0]=16'h0000;
		0707:	romdata[15:0]=16'h0000;
		0708:	romdata[15:0]=16'h0000;
		0709:	romdata[15:0]=16'h0000;
		0710:	romdata[15:0]=16'h0000;
		0711:	romdata[15:0]=16'h0000;
		0712:	romdata[15:0]=16'h0000;
		0713:	romdata[15:0]=16'h0000;
		0714:	romdata[15:0]=16'h0000;
		0715:	romdata[15:0]=16'h0000;
		0716:	romdata[15:0]=16'h0000;
		0717:	romdata[15:0]=16'h0000;
		0718:	romdata[15:0]=16'h0000;
		0719:	romdata[15:0]=16'h0000;
		0720:	romdata[15:0]=16'h0000;
		0721:	romdata[15:0]=16'h0000;
		0722:	romdata[15:0]=16'h0000;
		0723:	romdata[15:0]=16'h0000;
		0724:	romdata[15:0]=16'h0000;
		0725:	romdata[15:0]=16'h0000;
		0726:	romdata[15:0]=16'h0000;
		0727:	romdata[15:0]=16'h0000;
		0728:	romdata[15:0]=16'h0000;
		0729:	romdata[15:0]=16'h0000;
		0730:	romdata[15:0]=16'h0000;
		0731:	romdata[15:0]=16'h0000;
		0732:	romdata[15:0]=16'h0000;
		0733:	romdata[15:0]=16'h0000;
		0734:	romdata[15:0]=16'h0000;
		0735:	romdata[15:0]=16'h0000;
		0736:	romdata[15:0]=16'h0000;
		0737:	romdata[15:0]=16'h0000;
		0738:	romdata[15:0]=16'h0000;
		0739:	romdata[15:0]=16'h0000;
		0740:	romdata[15:0]=16'h0000;
		0741:	romdata[15:0]=16'h0000;
		0742:	romdata[15:0]=16'h0000;
		0743:	romdata[15:0]=16'h0000;
		0744:	romdata[15:0]=16'h0000;
		0745:	romdata[15:0]=16'h0000;
		0746:	romdata[15:0]=16'h0000;
		0747:	romdata[15:0]=16'h0000;
		0748:	romdata[15:0]=16'h0000;
		0749:	romdata[15:0]=16'h0000;
		0750:	romdata[15:0]=16'h0000;
		0751:	romdata[15:0]=16'h0000;
		0752:	romdata[15:0]=16'h0000;
		0753:	romdata[15:0]=16'h0000;
		0754:	romdata[15:0]=16'h0000;
		0755:	romdata[15:0]=16'h0000;
		0756:	romdata[15:0]=16'h0000;
		0757:	romdata[15:0]=16'h0000;
		0758:	romdata[15:0]=16'h0000;
		0759:	romdata[15:0]=16'h0000;
		0760:	romdata[15:0]=16'h0000;
		0761:	romdata[15:0]=16'h0000;
		0762:	romdata[15:0]=16'h0000;
		0763:	romdata[15:0]=16'h0000;
		0764:	romdata[15:0]=16'h0000;
		0765:	romdata[15:0]=16'h0000;
		0766:	romdata[15:0]=16'h0000;
		0767:	romdata[15:0]=16'h0000;
		0768:	romdata[15:0]=16'h0000;
		0769:	romdata[15:0]=16'h0000;
		0770:	romdata[15:0]=16'h0000;
		0771:	romdata[15:0]=16'h0000;
		0772:	romdata[15:0]=16'h0000;
		0773:	romdata[15:0]=16'h0000;
		0774:	romdata[15:0]=16'h0000;
		0775:	romdata[15:0]=16'h0000;
		0776:	romdata[15:0]=16'h0000;
		0777:	romdata[15:0]=16'h0000;
		0778:	romdata[15:0]=16'h0000;
		0779:	romdata[15:0]=16'h0000;
		0780:	romdata[15:0]=16'h0000;
		0781:	romdata[15:0]=16'h0000;
		0782:	romdata[15:0]=16'h0000;
		0783:	romdata[15:0]=16'h0000;
		0784:	romdata[15:0]=16'h0000;
		0785:	romdata[15:0]=16'h0000;
		0786:	romdata[15:0]=16'h0000;
		0787:	romdata[15:0]=16'h0000;
		0788:	romdata[15:0]=16'h0000;
		0789:	romdata[15:0]=16'h0000;
		0790:	romdata[15:0]=16'h0000;
		0791:	romdata[15:0]=16'h0000;
		0792:	romdata[15:0]=16'h0000;
		0793:	romdata[15:0]=16'h0000;
		0794:	romdata[15:0]=16'h0000;
		0795:	romdata[15:0]=16'h0000;
		0796:	romdata[15:0]=16'h0000;
		0797:	romdata[15:0]=16'h0000;
		0798:	romdata[15:0]=16'h0000;
		0799:	romdata[15:0]=16'h0000;
		0800:	romdata[15:0]=16'h0000;
		0801:	romdata[15:0]=16'h0000;
		0802:	romdata[15:0]=16'h0000;
		0803:	romdata[15:0]=16'h0000;
		0804:	romdata[15:0]=16'h0000;
		0805:	romdata[15:0]=16'h0000;
		0806:	romdata[15:0]=16'h0000;
		0807:	romdata[15:0]=16'h0000;
		0808:	romdata[15:0]=16'h0000;
		0809:	romdata[15:0]=16'h0000;
		0810:	romdata[15:0]=16'h0000;
		0811:	romdata[15:0]=16'h0000;
		0812:	romdata[15:0]=16'h0000;
		0813:	romdata[15:0]=16'h0000;
		0814:	romdata[15:0]=16'h0000;
		0815:	romdata[15:0]=16'h0000;
		0816:	romdata[15:0]=16'h0000;
		0817:	romdata[15:0]=16'h0000;
		0818:	romdata[15:0]=16'h0000;
		0819:	romdata[15:0]=16'h0000;
		0820:	romdata[15:0]=16'h0000;
		0821:	romdata[15:0]=16'h0000;
		0822:	romdata[15:0]=16'h0000;
		0823:	romdata[15:0]=16'h0000;
		0824:	romdata[15:0]=16'h0000;
		0825:	romdata[15:0]=16'h0000;
		0826:	romdata[15:0]=16'h0000;
		0827:	romdata[15:0]=16'h0000;
		0828:	romdata[15:0]=16'h0000;
		0829:	romdata[15:0]=16'h0000;
		0830:	romdata[15:0]=16'h0000;
		0831:	romdata[15:0]=16'h0000;
		0832:	romdata[15:0]=16'h0000;
		0833:	romdata[15:0]=16'h0000;
		0834:	romdata[15:0]=16'h0000;
		0835:	romdata[15:0]=16'h0000;
		0836:	romdata[15:0]=16'h0000;
		0837:	romdata[15:0]=16'h0000;
		0838:	romdata[15:0]=16'h0000;
		0839:	romdata[15:0]=16'h0000;
		0840:	romdata[15:0]=16'h0000;
		0841:	romdata[15:0]=16'h0000;
		0842:	romdata[15:0]=16'h0000;
		0843:	romdata[15:0]=16'h0000;
		0844:	romdata[15:0]=16'h0000;
		0845:	romdata[15:0]=16'h0000;
		0846:	romdata[15:0]=16'h0000;
		0847:	romdata[15:0]=16'h0000;
		0848:	romdata[15:0]=16'h0000;
		0849:	romdata[15:0]=16'h0000;
		0850:	romdata[15:0]=16'h0000;
		0851:	romdata[15:0]=16'h0000;
		0852:	romdata[15:0]=16'h0000;
		0853:	romdata[15:0]=16'h0000;
		0854:	romdata[15:0]=16'h0000;
		0855:	romdata[15:0]=16'h0000;
		0856:	romdata[15:0]=16'h0000;
		0857:	romdata[15:0]=16'h0000;
		0858:	romdata[15:0]=16'h0000;
		0859:	romdata[15:0]=16'h0000;
		0860:	romdata[15:0]=16'h0000;
		0861:	romdata[15:0]=16'h0000;
		0862:	romdata[15:0]=16'h0000;
		0863:	romdata[15:0]=16'h0000;
		0864:	romdata[15:0]=16'h0000;
		0865:	romdata[15:0]=16'h0000;
		0866:	romdata[15:0]=16'h0000;
		0867:	romdata[15:0]=16'h0000;
		0868:	romdata[15:0]=16'h0000;
		0869:	romdata[15:0]=16'h0000;
		0870:	romdata[15:0]=16'h0000;
		0871:	romdata[15:0]=16'h0000;
		0872:	romdata[15:0]=16'h0000;
		0873:	romdata[15:0]=16'h0000;
		0874:	romdata[15:0]=16'h0000;
		0875:	romdata[15:0]=16'h0000;
		0876:	romdata[15:0]=16'h0000;
		0877:	romdata[15:0]=16'h0000;
		0878:	romdata[15:0]=16'h0000;
		0879:	romdata[15:0]=16'h0000;
		0880:	romdata[15:0]=16'h0000;
		0881:	romdata[15:0]=16'h0000;
		0882:	romdata[15:0]=16'h0000;
		0883:	romdata[15:0]=16'h0000;
		0884:	romdata[15:0]=16'h0000;
		0885:	romdata[15:0]=16'h0000;
		0886:	romdata[15:0]=16'h0000;
		0887:	romdata[15:0]=16'h0000;
		0888:	romdata[15:0]=16'h0000;
		0889:	romdata[15:0]=16'h0000;
		0890:	romdata[15:0]=16'h0000;
		0891:	romdata[15:0]=16'h0000;
		0892:	romdata[15:0]=16'h0000;
		0893:	romdata[15:0]=16'h0000;
		0894:	romdata[15:0]=16'h0000;
		0895:	romdata[15:0]=16'h0000;
		0896:	romdata[15:0]=16'h0000;
		0897:	romdata[15:0]=16'h0000;
		0898:	romdata[15:0]=16'h0000;
		0899:	romdata[15:0]=16'h0000;
		0900:	romdata[15:0]=16'h0000;
		0901:	romdata[15:0]=16'h0000;
		0902:	romdata[15:0]=16'h0000;
		0903:	romdata[15:0]=16'h0000;
		0904:	romdata[15:0]=16'h0000;
		0905:	romdata[15:0]=16'h0000;
		0906:	romdata[15:0]=16'h0000;
		0907:	romdata[15:0]=16'h0000;
		0908:	romdata[15:0]=16'h0000;
		0909:	romdata[15:0]=16'h0000;
		0910:	romdata[15:0]=16'h0000;
		0911:	romdata[15:0]=16'h0000;
		0912:	romdata[15:0]=16'h0000;
		0913:	romdata[15:0]=16'h0000;
		0914:	romdata[15:0]=16'h0000;
		0915:	romdata[15:0]=16'h0000;
		0916:	romdata[15:0]=16'h0000;
		0917:	romdata[15:0]=16'h0000;
		0918:	romdata[15:0]=16'h0000;
		0919:	romdata[15:0]=16'h0000;
		0920:	romdata[15:0]=16'h0000;
		0921:	romdata[15:0]=16'h0000;
		0922:	romdata[15:0]=16'h0000;
		0923:	romdata[15:0]=16'h0000;
		0924:	romdata[15:0]=16'h0000;
		0925:	romdata[15:0]=16'h0000;
		0926:	romdata[15:0]=16'h0000;
		0927:	romdata[15:0]=16'h0000;
		0928:	romdata[15:0]=16'h0000;
		0929:	romdata[15:0]=16'h0000;
		0930:	romdata[15:0]=16'h0000;
		0931:	romdata[15:0]=16'h0000;
		0932:	romdata[15:0]=16'h0000;
		0933:	romdata[15:0]=16'h0000;
		0934:	romdata[15:0]=16'h0000;
		0935:	romdata[15:0]=16'h0000;
		0936:	romdata[15:0]=16'h0000;
		0937:	romdata[15:0]=16'h0000;
		0938:	romdata[15:0]=16'h0000;
		0939:	romdata[15:0]=16'h0000;
		0940:	romdata[15:0]=16'h0000;
		0941:	romdata[15:0]=16'h0000;
		0942:	romdata[15:0]=16'h0000;
		0943:	romdata[15:0]=16'h0000;
		0944:	romdata[15:0]=16'h0000;
		0945:	romdata[15:0]=16'h0000;
		0946:	romdata[15:0]=16'h0000;
		0947:	romdata[15:0]=16'h0000;
		0948:	romdata[15:0]=16'h0000;
		0949:	romdata[15:0]=16'h0000;
		0950:	romdata[15:0]=16'h0000;
		0951:	romdata[15:0]=16'h0000;
		0952:	romdata[15:0]=16'h0000;
		0953:	romdata[15:0]=16'h0000;
		0954:	romdata[15:0]=16'h0000;
		0955:	romdata[15:0]=16'h0000;
		0956:	romdata[15:0]=16'h0000;
		0957:	romdata[15:0]=16'h0000;
		0958:	romdata[15:0]=16'h0000;
		0959:	romdata[15:0]=16'h0000;
		0960:	romdata[15:0]=16'h0000;
		0961:	romdata[15:0]=16'h0000;
		0962:	romdata[15:0]=16'h0000;
		0963:	romdata[15:0]=16'h0000;
		0964:	romdata[15:0]=16'h0000;
		0965:	romdata[15:0]=16'h0000;
		0966:	romdata[15:0]=16'h0000;
		0967:	romdata[15:0]=16'h0000;
		0968:	romdata[15:0]=16'h0000;
		0969:	romdata[15:0]=16'h0000;
		0970:	romdata[15:0]=16'h0000;
		0971:	romdata[15:0]=16'h0000;
		0972:	romdata[15:0]=16'h0000;
		0973:	romdata[15:0]=16'h0000;
		0974:	romdata[15:0]=16'h0000;
		0975:	romdata[15:0]=16'h0000;
		0976:	romdata[15:0]=16'h0000;
		0977:	romdata[15:0]=16'h0000;
		0978:	romdata[15:0]=16'h0000;
		0979:	romdata[15:0]=16'h0000;
		0980:	romdata[15:0]=16'h0000;
		0981:	romdata[15:0]=16'h0000;
		0982:	romdata[15:0]=16'h0000;
		0983:	romdata[15:0]=16'h0000;
		0984:	romdata[15:0]=16'h0000;
		0985:	romdata[15:0]=16'h0000;
		0986:	romdata[15:0]=16'h0000;
		0987:	romdata[15:0]=16'h0000;
		0988:	romdata[15:0]=16'h0000;
		0989:	romdata[15:0]=16'h0000;
		0990:	romdata[15:0]=16'h0000;
		0991:	romdata[15:0]=16'h0000;
		0992:	romdata[15:0]=16'h0000;
		0993:	romdata[15:0]=16'h0000;
		0994:	romdata[15:0]=16'h0000;
		0995:	romdata[15:0]=16'h0000;
		0996:	romdata[15:0]=16'h0000;
		0997:	romdata[15:0]=16'h0000;
		0998:	romdata[15:0]=16'h0000;
		0999:	romdata[15:0]=16'h0000;
		1000:	romdata[15:0]=16'h0000;
		1001:	romdata[15:0]=16'h0000;
		1002:	romdata[15:0]=16'h0000;
		1003:	romdata[15:0]=16'h0000;
		1004:	romdata[15:0]=16'h0000;
		1005:	romdata[15:0]=16'h0000;
		1006:	romdata[15:0]=16'h0000;
		1007:	romdata[15:0]=16'h0000;
		1008:	romdata[15:0]=16'h0000;
		1009:	romdata[15:0]=16'h0000;
		1010:	romdata[15:0]=16'h0000;
		1011:	romdata[15:0]=16'h0000;
		1012:	romdata[15:0]=16'h0000;
		1013:	romdata[15:0]=16'h0000;
		1014:	romdata[15:0]=16'h0000;
		1015:	romdata[15:0]=16'h0000;
		1016:	romdata[15:0]=16'h0000;
		1017:	romdata[15:0]=16'h0000;
		1018:	romdata[15:0]=16'h0000;
		1019:	romdata[15:0]=16'h0000;
		1020:	romdata[15:0]=16'h0000;
		1021:	romdata[15:0]=16'h0000;
		1022:	romdata[15:0]=16'h0000;
		1023:	romdata[15:0]=16'h0000;
	endcase
end

 //output enable
always @(romdata or aen or rd)
	if(aen && rd)
		dataout[15:0]=romdata[15:0];
	else
		dataout[15:0]=16'h0000;

endmodule
